`default_nettype none
`timescale 1ns / 1ps

module top(
    input wire clk,
    input wire btnc,
);

endmodule
